magic
tech sky130A
magscale 1 2
timestamp 1605225592
<< nwell >>
rect -300 309 300 630
<< nmos >>
rect -180 90 -150 180
rect -70 90 -40 180
rect 40 90 70 180
rect 150 90 180 180
<< pmos >>
rect -180 460 -150 550
rect -70 460 -40 550
rect 40 460 70 550
rect 150 460 180 550
<< ndiff >>
rect -260 160 -180 180
rect -260 120 -240 160
rect -200 120 -180 160
rect -260 90 -180 120
rect -150 170 -70 180
rect -150 130 -130 170
rect -90 130 -70 170
rect -150 90 -70 130
rect -40 150 40 180
rect -40 110 -20 150
rect 20 110 40 150
rect -40 90 40 110
rect 70 170 150 180
rect 70 130 90 170
rect 130 130 150 170
rect 70 90 150 130
rect 180 160 260 180
rect 180 120 200 160
rect 240 120 260 160
rect 180 90 260 120
<< pdiff >>
rect -260 520 -180 550
rect -260 480 -240 520
rect -200 480 -180 520
rect -260 460 -180 480
rect -150 460 -70 550
rect -40 530 40 550
rect -40 490 -20 530
rect 20 490 40 530
rect -40 460 40 490
rect 70 460 150 550
rect 180 520 260 550
rect 180 480 200 520
rect 240 480 260 520
rect 180 460 260 480
<< ndiffc >>
rect -240 120 -200 160
rect -130 130 -90 170
rect -20 110 20 150
rect 90 130 130 170
rect 200 120 240 160
<< pdiffc >>
rect -240 480 -200 520
rect -20 490 20 530
rect 200 480 240 520
<< poly >>
rect -180 550 -150 580
rect -70 550 -40 580
rect 40 550 70 580
rect 150 550 180 580
rect -180 410 -150 460
rect -240 390 -150 410
rect -240 350 -230 390
rect -190 350 -150 390
rect -70 380 -40 460
rect -240 330 -150 350
rect -180 180 -150 330
rect -76 370 -4 380
rect -76 330 -60 370
rect -20 330 -4 370
rect -76 320 -4 330
rect -70 180 -40 320
rect 40 270 70 460
rect 150 410 180 460
rect 150 390 240 410
rect 150 350 190 390
rect 230 350 240 390
rect 150 330 240 350
rect 4 260 76 270
rect 4 220 20 260
rect 60 220 76 260
rect 4 210 76 220
rect 40 180 70 210
rect 150 180 180 330
rect -180 60 -150 90
rect -70 60 -40 90
rect 40 60 70 90
rect 150 60 180 90
<< polycont >>
rect -230 350 -190 390
rect -60 330 -20 370
rect 190 350 230 390
rect 20 220 60 260
<< locali >>
rect -150 606 -130 610
rect -260 572 -130 606
rect -150 570 -130 572
rect -90 570 -20 610
rect 20 570 90 610
rect 130 606 150 610
rect 130 572 260 606
rect 130 570 150 572
rect -20 530 20 570
rect -256 480 -240 520
rect -200 480 -110 520
rect -230 390 -190 410
rect -230 330 -190 350
rect -150 280 -110 480
rect -20 470 20 490
rect 80 480 200 520
rect 240 480 256 520
rect -76 370 -4 380
rect 80 370 120 480
rect 190 390 230 410
rect -76 330 -60 370
rect -20 330 150 370
rect 190 330 230 350
rect -76 320 -4 330
rect -150 270 40 280
rect -150 260 76 270
rect -150 240 20 260
rect -240 160 -200 220
rect -240 100 -200 120
rect -130 170 -90 240
rect 0 220 20 240
rect 60 220 76 260
rect 0 210 76 220
rect 110 170 150 330
rect -130 110 -90 130
rect -20 150 20 170
rect 74 130 90 170
rect 130 130 150 170
rect 200 160 240 220
rect -20 70 20 110
rect 200 100 240 120
rect -150 65 -130 70
rect -260 31 -130 65
rect -150 30 -130 31
rect -90 30 -20 70
rect 20 30 90 70
rect 130 65 150 70
rect 130 31 260 65
rect 130 30 150 31
<< viali >>
rect -130 570 -90 610
rect -20 570 20 610
rect 90 570 130 610
rect -230 350 -190 390
rect 190 350 230 390
rect -130 30 -90 70
rect -20 30 20 70
rect 90 30 130 70
<< metal1 >>
rect -260 610 260 640
rect -260 570 -130 610
rect -90 570 -20 610
rect 20 570 90 610
rect 130 570 260 610
rect -260 544 260 570
rect -220 430 220 470
rect -220 410 -180 430
rect -240 390 -180 410
rect -240 350 -230 390
rect -190 350 -180 390
rect -240 330 -180 350
rect 180 410 220 430
rect 180 390 240 410
rect 180 350 190 390
rect 230 350 240 390
rect 180 330 240 350
rect -260 70 260 96
rect -260 30 -130 70
rect -90 30 -20 70
rect 20 30 90 70
rect 130 30 260 70
rect -260 0 260 30
<< labels >>
rlabel metal1 180 330 240 410 0 EN
rlabel metal1 -240 330 -180 410 0 EN
rlabel locali 20 220 60 260 0 Q
rlabel locali -60 330 -20 370 0 Q_N
rlabel locali 200 180 240 220 0 D_N
rlabel locali -240 180 -200 220 0 D
rlabel nwell -300 309 300 630 1 NWELL
rlabel viali -20 570 20 610 1 VPWR
rlabel viali -20 30 20 70 1 VGND
<< end >>
