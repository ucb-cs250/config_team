DLatch Simulation

.lib "./sky130_fd_pr/models/sky130.lib.spice" tt 

Vgnd VGND 0 0
Vdd VPWR VGND 1.8

Ven EN  VGND pulse(0 1.8 0.5n  10p 10p 1n 2n)

Vd  D   VGND pulse(0 1.8 3.75n 10p 10p 5n 10n)
vdn D_N VGND pulse(1.8 0 3.75n 10p 10p 5n 10n)

// R1 Q VPWR 100k
// R2 Q_N VPWR 100k

.tran 10e-12 10e-09 0e-00

.control
run
plot EN D D_N Q Q_N
.endc

.subckt dlatchp EN D D_N Q Q_N VGND VPWR NWELL VSUBS
X0 a_n150_460# EN Q NWELL sky130_fd_pr__pfet_01v8 w=450000u l=150000u
X1 D_N EN Q_N VSUBS sky130_fd_pr__nfet_01v8 w=450000u l=150000u
X2 Q_N EN a_70_460# NWELL sky130_fd_pr__pfet_01v8 w=450000u l=150000u
X3 a_70_460# Q VPWR NWELL sky130_fd_pr__pfet_01v8 w=450000u l=150000u
X4 Q_N Q VGND VSUBS sky130_fd_pr__nfet_01v8 w=450000u l=150000u
X5 VPWR Q_N a_n150_460# NWELL sky130_fd_pr__pfet_01v8 w=450000u l=150000u
X6 Q EN D VSUBS sky130_fd_pr__nfet_01v8 w=450000u l=150000u
X7 VGND Q_N Q VSUBS sky130_fd_pr__nfet_01v8 w=450000u l=150000u
C0 D Q_N 0.01fF
C1 VPWR D_N 0.00fF
C2 Q_N NWELL 0.01fF
C3 D VGND 0.07fF
C4 D_N Q_N 0.06fF
C5 a_70_460# EN 0.02fF
C6 a_n150_460# EN 0.02fF
C7 D_N VGND 0.07fF
C8 a_n150_460# Q 0.03fF
C9 a_70_460# VPWR 0.02fF
C10 a_n150_460# VPWR 0.02fF
C11 a_70_460# Q_N 0.05fF
C12 EN Q 0.42fF
C13 VPWR EN 0.39fF
C14 VPWR Q 0.18fF
C15 EN Q_N 0.41fF
C16 EN VGND 0.14fF
C17 Q_N Q 0.47fF
C18 EN D 0.01fF
C19 VPWR Q_N 0.23fF
C20 VGND Q 0.16fF
C21 EN NWELL 0.01fF
C22 D Q 0.06fF
C23 EN D_N 0.01fF
C24 VPWR VGND 0.00fF
C25 VPWR D 0.00fF
C26 Q NWELL 0.01fF
C27 D_N Q 0.02fF
C28 VPWR NWELL 0.03fF
C29 VGND Q_N 0.14fF
C30 D_N VSUBS 0.03fF
C31 VGND VSUBS 0.42fF
C32 D VSUBS 0.03fF
C33 VPWR VSUBS 0.41fF
C34 Q VSUBS 0.45fF
C35 Q_N VSUBS 0.45fF
C36 EN VSUBS 0.69fF
C37 NWELL VSUBS 0.58fF
.ends


Xdlatchpinst EN D D_N Q Q_N VGND VPWR NWELL VSUBS dlatchp

.end
