magic
tech sky130A
magscale 1 2
timestamp 1605251239
<< nwell >>
rect -300 309 300 630
<< nmos >>
rect -180 90 -150 180
rect -70 90 -40 180
rect 40 90 70 180
rect 150 90 180 180
<< pmos >>
rect -180 460 -150 550
rect -70 460 -40 550
rect 40 460 70 550
rect 150 460 180 550
<< ndiff >>
rect -260 150 -180 180
rect -260 110 -240 150
rect -200 110 -180 150
rect -260 90 -180 110
rect -150 90 -70 180
rect -40 150 40 180
rect -40 110 -20 150
rect 20 110 40 150
rect -40 90 40 110
rect 70 90 150 180
rect 180 150 260 180
rect 180 110 200 150
rect 240 110 260 150
rect 180 90 260 110
<< pdiff >>
rect -260 520 -180 550
rect -260 480 -240 520
rect -200 480 -180 520
rect -260 460 -180 480
rect -150 510 -70 550
rect -150 470 -130 510
rect -90 470 -70 510
rect -150 460 -70 470
rect -40 530 40 550
rect -40 490 -20 530
rect 20 490 40 530
rect -40 460 40 490
rect 70 510 150 550
rect 70 470 90 510
rect 130 470 150 510
rect 70 460 150 470
rect 180 520 260 550
rect 180 480 200 520
rect 240 480 260 520
rect 180 460 260 480
<< ndiffc >>
rect -240 110 -200 150
rect -20 110 20 150
rect 200 110 240 150
<< pdiffc >>
rect -240 480 -200 520
rect -130 470 -90 510
rect -20 490 20 530
rect 90 470 130 510
rect 200 480 240 520
<< poly >>
rect -180 550 -150 580
rect -70 550 -40 580
rect 40 550 70 580
rect 150 550 180 580
rect -180 310 -150 460
rect -240 290 -150 310
rect -240 250 -230 290
rect -190 250 -150 290
rect -70 270 -40 460
rect 40 380 70 460
rect 4 370 76 380
rect 4 330 20 370
rect 60 330 76 370
rect 4 320 76 330
rect -240 230 -150 250
rect -180 180 -150 230
rect -76 260 -4 270
rect -76 220 -60 260
rect -20 220 -4 260
rect -76 210 -4 220
rect -70 180 -40 210
rect 40 180 70 320
rect 150 310 180 460
rect 150 290 240 310
rect 150 250 190 290
rect 230 250 240 290
rect 150 230 240 250
rect 150 180 180 230
rect -180 60 -150 90
rect -70 60 -40 90
rect 40 60 70 90
rect 150 60 180 90
<< polycont >>
rect -230 250 -190 290
rect 20 330 60 370
rect -60 220 -20 260
rect 190 250 230 290
<< locali >>
rect -150 606 -130 610
rect -260 572 -130 606
rect -150 570 -130 572
rect -90 570 -20 610
rect 20 570 90 610
rect 130 606 150 610
rect 130 572 260 606
rect 130 570 150 572
rect -240 520 -200 536
rect -20 530 20 570
rect -240 420 -200 480
rect -150 470 -130 510
rect -90 470 -70 510
rect 200 520 240 536
rect -20 470 20 490
rect 70 470 90 510
rect 130 470 150 510
rect -150 370 -110 470
rect 4 370 76 380
rect -150 330 20 370
rect 60 330 76 370
rect -230 290 -190 310
rect -230 230 -190 250
rect -150 150 -110 330
rect 4 320 76 330
rect -76 260 -4 270
rect 110 260 150 470
rect 200 420 240 480
rect -76 220 -60 260
rect -20 220 150 260
rect 190 290 230 310
rect 190 230 230 250
rect -76 210 -4 220
rect -256 110 -240 150
rect -200 110 -110 150
rect -20 150 20 170
rect 110 150 150 220
rect 110 110 200 150
rect 240 110 256 150
rect -20 70 20 110
rect -150 65 -130 70
rect -260 31 -130 65
rect -150 30 -130 31
rect -90 30 -20 70
rect 20 30 90 70
rect 130 65 150 70
rect 130 31 260 65
rect 130 30 150 31
<< viali >>
rect -130 570 -90 610
rect -20 570 20 610
rect 90 570 130 610
rect -230 250 -190 290
rect 190 250 230 290
rect -130 30 -90 70
rect -20 30 20 70
rect 90 30 130 70
<< metal1 >>
rect -260 610 260 640
rect -260 570 -130 610
rect -90 570 -20 610
rect 20 570 90 610
rect 130 570 260 610
rect -260 544 260 570
rect -240 290 -180 310
rect -240 250 -230 290
rect -190 250 -180 290
rect -240 230 -180 250
rect -220 210 -180 230
rect 180 290 240 310
rect 180 250 190 290
rect 230 250 240 290
rect 180 230 240 250
rect 180 210 220 230
rect -220 170 220 210
rect -260 70 260 96
rect -260 30 -130 70
rect -90 30 -20 70
rect 20 30 90 70
rect 130 30 260 70
rect -260 0 260 30
<< labels >>
rlabel nwell -300 309 300 630 1 NWELL
rlabel viali -20 570 20 610 1 VPWR
rlabel viali -20 30 20 70 1 VGND
rlabel locali 20 330 60 370 0 Q_N
rlabel locali -60 220 -20 260 0 Q
rlabel metal1 -240 230 -180 310 0 EN
rlabel metal1 180 230 240 310 0 EN
rlabel locali -240 420 -200 460 0 D_N
rlabel locali 200 420 240 460 0 D
<< end >>
