`timescale 1ns/1ps

`include "../behavioral/config_sram_data.v"

module config_sram_data_tb_top;
    initial begin
    end
endmodule // config_sram_data_tb_top
