`timescale 1ns/1ps

`include "../behavioral/config_tile.v"

module config_tile_tb_top;
    initial begin
    end
endmodule // config_tile_tb_top
